﻿// TB: simulate PTEST/PFLUSH/PLOAD/MOVEC sequences
