﻿// TB: TLB hit/miss/refill + PFLUSH
