﻿// TB: perms
