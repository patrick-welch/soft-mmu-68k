﻿// TB: descriptor pack/unpack
