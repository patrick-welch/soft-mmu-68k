﻿// checkers, scoreboards (sim-only)
