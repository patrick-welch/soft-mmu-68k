﻿// typedefs/structs (sim-only)
