﻿// TB: VAâ†’PA + faults + TTR bypass
