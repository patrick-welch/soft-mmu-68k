﻿// TB: walker
